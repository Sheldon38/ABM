module bus #(parameter WIDTH=8)(
inout wire [WIDTH-1:0] datapath
);
endmodule